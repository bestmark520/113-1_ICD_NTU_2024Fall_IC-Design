* SPICE NETLIST
***************************************

*.CALIBRE ABORT_INFO SOFTCHK
.SUBCKT L POS NEG
.ENDS
***************************************
.SUBCKT inv3 1 2 3
** N=5 EP=3 IP=0 FDC=2

*M0 4 1 3 3 N
M0 4 1 2 3 N_18 L=1.8e-07 W=2e-06 AD=1.52e-12 AS=1.8e-12 PD=3.52e-06 PS=3.8e-06 $X=1400 $Y=-2680 $D=0
M1 4 1 5 5 P_18 L=1.8e-07 W=2.5e-06 AD=1.9e-12 AS=2.25e-12 PD=4.02e-06 PS=4.3e-06 $X=1400 $Y=1000 $D=1
.ENDS
***************************************
.SUBCKT n_mos_GND 1 2 3 4
** N=4 EP=4 IP=0 FDC=1
M0 1 2 3 4 N_18 L=1.8e-07 W=2e-06 AD=1.52e-12 AS=1.8e-12 PD=3.52e-06 PS=3.8e-06 $X=1400 $Y=-2680 $D=0
.ENDS
***************************************
.SUBCKT p_mos 1 2 3
** N=5 EP=3 IP=0 FDC=1
M0 1 3 2 5 P_18 L=1.8e-07 W=2.5e-06 AD=1.9e-12 AS=2.25e-12 PD=4.02e-06 PS=4.3e-06 $X=1400 $Y=1000 $D=1
.ENDS
***************************************
.SUBCKT n_mos 1 2 3 5
** N=5 EP=4 IP=0 FDC=1
M0 1 3 2 5 N_18 L=1.8e-07 W=2e-06 AD=1.52e-12 AS=1.8e-12 PD=3.52e-06 PS=3.8e-06 $X=1400 $Y=-2680 $D=0
.ENDS
***************************************
.SUBCKT p_mos_VDD 1 2
** N=4 EP=2 IP=0 FDC=1
M0 1 2 4 4 P_18 L=1.8e-07 W=2.5e-06 AD=1.9e-12 AS=2.25e-12 PD=4.02e-06 PS=4.3e-06 $X=1400 $Y=1000 $D=1
.ENDS
***************************************
.SUBCKT adder
** N=31 EP=0 IP=100 FDC=28
X0 5 18 18 inv3 $T=-25350 -18680 0 0 $X=-26550 $Y=-23960
X1 11 19 18 inv3 $T=85340 2750 0 0 $X=84140 $Y=-2530
X2 1 12 20 18 n_mos_GND $T=-70190 -1710 0 0 $X=-70790 $Y=-6990
X3 1 4 21 18 n_mos_GND $T=-55430 -1710 0 0 $X=-56030 $Y=-6990
X4 4 4 22 18 n_mos_GND $T=-7110 27390 0 0 $X=-7710 $Y=22110
X5 8 12 23 18 n_mos_GND $T=-5990 -1710 0 0 $X=-6590 $Y=-6990
X6 8 4 24 18 n_mos_GND $T=32390 -1710 0 0 $X=31790 $Y=-6990
X7 8 13 25 18 n_mos_GND $T=45890 -1710 0 0 $X=45290 $Y=-6990
X8 10 13 26 18 n_mos_GND $T=66810 27390 0 0 $X=66210 $Y=22110
X9 2 14 13 p_mos $T=-40250 8970 0 0 $X=-41750 $Y=8360
X10 5 3 4 p_mos $T=-5500 34680 0 0 $X=-7000 $Y=34070
X11 11 5 8 p_mos $T=11630 8530 0 0 $X=10130 $Y=7920
X12 9 15 4 p_mos $T=50520 34680 0 0 $X=49020 $Y=34070
X13 11 16 13 p_mos $T=66210 34680 0 0 $X=64710 $Y=34070
X14 1 17 13 18 n_mos $T=-40340 -1810 0 0 $X=-41540 $Y=-7090
X15 5 4 12 18 n_mos $T=-19840 27380 0 0 $X=-21040 $Y=22100
X16 11 5 8 18 n_mos $T=11470 -1810 0 0 $X=10270 $Y=-7090
X17 11 7 12 18 n_mos $T=33570 27380 0 0 $X=32370 $Y=22100
X18 7 10 4 18 n_mos $T=50950 27380 0 0 $X=49750 $Y=22100
X19 2 12 p_mos_VDD $T=-69940 8470 0 0 $X=-71140 $Y=7860
X20 2 4 p_mos_VDD $T=-55100 8470 0 0 $X=-56300 $Y=7860
X21 3 12 p_mos_VDD $T=-20080 34270 0 0 $X=-21280 $Y=33660
X22 8 12 p_mos_VDD $T=-5730 8030 0 0 $X=-6930 $Y=7420
X23 8 4 p_mos_VDD $T=32660 8030 0 0 $X=31460 $Y=7420
X24 6 12 p_mos_VDD $T=33580 34270 0 0 $X=32380 $Y=33660
X25 8 13 p_mos_VDD $T=45910 8030 0 0 $X=44710 $Y=7420
*.CALIBRE WARNING SCONNECT SCONNECT conflict(s) detected by extraction in this cell. See extraction report for details.
.ENDS
***************************************
