* SPICE NETLIST
***************************************

.SUBCKT L POS NEG
.ENDS
***************************************
.SUBCKT n_mos GND
** N=4 EP=1 IP=0 FDC=1
M0 1 3 2 GND N_18 L=1.8e-07 W=2e-06 AD=1.52e-12 AS=1.8e-12 PD=3.52e-06 PS=3.8e-06 $X=1400 $Y=-2680 $D=0
.ENDS
***************************************
