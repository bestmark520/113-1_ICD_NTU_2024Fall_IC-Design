* SPICE NETLIST
***************************************

.SUBCKT L POS NEG
.ENDS
***************************************
.SUBCKT inv3 1 2 3 4
** N=4 EP=4 IP=0 FDC=2
M0 1 2 3 3 N_18 L=1.8e-07 W=2e-06 AD=1.52e-12 AS=1.8e-12 PD=3.52e-06 PS=3.8e-06 $X=1400 $Y=-2680 $D=0
M1 1 2 4 4 P_18 L=1.8e-07 W=2.5e-06 AD=1.9e-12 AS=2.25e-12 PD=4.02e-06 PS=4.3e-06 $X=1400 $Y=1000 $D=1
.ENDS
***************************************
.SUBCKT n_mos_GND 1 2 3
** N=3 EP=3 IP=0 FDC=1
M0 1 2 3 3 N_18 L=1.8e-07 W=2e-06 AD=1.52e-12 AS=1.8e-12 PD=3.52e-06 PS=3.8e-06 $X=1400 $Y=-2680 $D=0
.ENDS
***************************************
.SUBCKT p_mos 1 2 3 4
** N=5 EP=4 IP=0 FDC=1
M0 1 3 2 4 P_18 L=1.8e-07 W=2.5e-06 AD=1.9e-12 AS=2.25e-12 PD=4.02e-06 PS=4.3e-06 $X=1400 $Y=1000 $D=1
.ENDS
***************************************
.SUBCKT n_mos 1 2 3 4
** N=4 EP=4 IP=0 FDC=1
M0 1 3 2 4 N_18 L=1.8e-07 W=2e-06 AD=1.52e-12 AS=1.8e-12 PD=3.52e-06 PS=3.8e-06 $X=1400 $Y=-2680 $D=0
.ENDS
***************************************
.SUBCKT p_mos_VDD 1 2 3
** N=4 EP=3 IP=0 FDC=1
M0 1 2 3 3 P_18 L=1.8e-07 W=2.5e-06 AD=1.9e-12 AS=2.25e-12 PD=4.02e-06 PS=4.3e-06 $X=1400 $Y=1000 $D=1
.ENDS
***************************************
.SUBCKT adder C1 C2 C3 S1 S2 S3 Cout S4 A1 B1 Cin A2 B2 A3 B3 A4 B4 GND VDD
** N=67 EP=19 IP=408 FDC=112
X0 C1 5 GND VDD inv3 $T=-25180 -18620 0 0 $X=-26380 $Y=-23900
X1 S1 12 GND VDD inv3 $T=84940 2760 0 0 $X=83740 $Y=-2520
X2 C2 18 GND VDD inv3 $T=143450 -18620 0 0 $X=142250 $Y=-23900
X3 S2 25 GND VDD inv3 $T=253570 2760 0 0 $X=252370 $Y=-2520
X4 C3 31 GND VDD inv3 $T=311320 -18620 0 0 $X=310120 $Y=-23900
X5 S3 38 GND VDD inv3 $T=421020 2760 0 0 $X=419820 $Y=-2520
X6 Cout 44 GND VDD inv3 $T=481470 -18620 0 0 $X=480270 $Y=-23900
X7 S4 51 GND VDD inv3 $T=591590 2760 0 0 $X=590390 $Y=-2520
X8 2 A1 GND n_mos_GND $T=-70190 -1710 0 0 $X=-70790 $Y=-6990
X9 2 B1 GND n_mos_GND $T=-55430 -1710 0 0 $X=-56030 $Y=-6990
X10 4 B1 GND n_mos_GND $T=-7110 27390 0 0 $X=-7710 $Y=22110
X11 7 A1 GND n_mos_GND $T=-5990 -1710 0 0 $X=-6590 $Y=-6990
X12 7 B1 GND n_mos_GND $T=32390 -1710 0 0 $X=31790 $Y=-6990
X13 7 Cin GND n_mos_GND $T=45890 -1710 0 0 $X=45290 $Y=-6990
X14 11 Cin GND n_mos_GND $T=66810 27390 0 0 $X=66210 $Y=22110
X15 15 A2 GND n_mos_GND $T=98440 -1710 0 0 $X=97840 $Y=-6990
X16 15 B2 GND n_mos_GND $T=113200 -1710 0 0 $X=112600 $Y=-6990
X17 17 B2 GND n_mos_GND $T=161520 27390 0 0 $X=160920 $Y=22110
X18 20 A2 GND n_mos_GND $T=162640 -1710 0 0 $X=162040 $Y=-6990
X19 20 B2 GND n_mos_GND $T=201020 -1710 0 0 $X=200420 $Y=-6990
X20 20 C1 GND n_mos_GND $T=214520 -1710 0 0 $X=213920 $Y=-6990
X21 24 C1 GND n_mos_GND $T=235440 27390 0 0 $X=234840 $Y=22110
X22 28 A3 GND n_mos_GND $T=266310 -1710 0 0 $X=265710 $Y=-6990
X23 28 B3 GND n_mos_GND $T=281070 -1710 0 0 $X=280470 $Y=-6990
X24 30 B3 GND n_mos_GND $T=329390 27390 0 0 $X=328790 $Y=22110
X25 33 A3 GND n_mos_GND $T=330510 -1710 0 0 $X=329910 $Y=-6990
X26 33 B3 GND n_mos_GND $T=368890 -1710 0 0 $X=368290 $Y=-6990
X27 33 C2 GND n_mos_GND $T=382390 -1710 0 0 $X=381790 $Y=-6990
X28 37 C2 GND n_mos_GND $T=403310 27390 0 0 $X=402710 $Y=22110
X29 41 A4 GND n_mos_GND $T=436460 -1710 0 0 $X=435860 $Y=-6990
X30 41 B4 GND n_mos_GND $T=451220 -1710 0 0 $X=450620 $Y=-6990
X31 43 B4 GND n_mos_GND $T=499540 27390 0 0 $X=498940 $Y=22110
X32 46 A4 GND n_mos_GND $T=500660 -1710 0 0 $X=500060 $Y=-6990
X33 46 B4 GND n_mos_GND $T=539040 -1710 0 0 $X=538440 $Y=-6990
X34 46 C3 GND n_mos_GND $T=552540 -1710 0 0 $X=551940 $Y=-6990
X35 50 C3 GND n_mos_GND $T=573460 27390 0 0 $X=572860 $Y=22110
X36 5 1 Cin VDD p_mos $T=-40250 8970 0 0 $X=-41750 $Y=8360
X37 5 3 B1 VDD p_mos $T=-5500 34680 0 0 $X=-7000 $Y=34070
X38 12 9 5 VDD p_mos $T=11630 8530 0 0 $X=10130 $Y=7920
X39 10 6 B1 VDD p_mos $T=50520 34680 0 0 $X=49020 $Y=34070
X40 12 10 Cin VDD p_mos $T=66210 34680 0 0 $X=64710 $Y=34070
X41 18 14 C1 VDD p_mos $T=128380 8970 0 0 $X=126880 $Y=8360
X42 18 16 B2 VDD p_mos $T=163130 34680 0 0 $X=161630 $Y=34070
X43 25 22 18 VDD p_mos $T=180260 8530 0 0 $X=178760 $Y=7920
X44 23 19 B2 VDD p_mos $T=219150 34680 0 0 $X=217650 $Y=34070
X45 25 23 C1 VDD p_mos $T=234840 34680 0 0 $X=233340 $Y=34070
X46 31 27 C2 VDD p_mos $T=296250 8970 0 0 $X=294750 $Y=8360
X47 31 29 B3 VDD p_mos $T=331000 34680 0 0 $X=329500 $Y=34070
X48 38 35 31 VDD p_mos $T=348130 8530 0 0 $X=346630 $Y=7920
X49 36 32 B3 VDD p_mos $T=387020 34680 0 0 $X=385520 $Y=34070
X50 38 36 C2 VDD p_mos $T=402710 34680 0 0 $X=401210 $Y=34070
X51 44 40 C3 VDD p_mos $T=466400 8970 0 0 $X=464900 $Y=8360
X52 44 42 B4 VDD p_mos $T=501150 34680 0 0 $X=499650 $Y=34070
X53 51 48 44 VDD p_mos $T=518280 8530 0 0 $X=516780 $Y=7920
X54 49 45 B4 VDD p_mos $T=557170 34680 0 0 $X=555670 $Y=34070
X55 51 49 C3 VDD p_mos $T=572860 34680 0 0 $X=571360 $Y=34070
X56 5 2 Cin GND n_mos $T=-40340 -1810 0 0 $X=-41540 $Y=-7090
X57 5 4 A1 GND n_mos $T=-19840 27380 0 0 $X=-21040 $Y=22100
X58 12 7 5 GND n_mos $T=11470 -1810 0 0 $X=10270 $Y=-7090
X59 12 8 A1 GND n_mos $T=33570 27380 0 0 $X=32370 $Y=22100
X60 8 11 B1 GND n_mos $T=50950 27380 0 0 $X=49750 $Y=22100
X61 18 15 C1 GND n_mos $T=128290 -1810 0 0 $X=127090 $Y=-7090
X62 18 17 A2 GND n_mos $T=148790 27380 0 0 $X=147590 $Y=22100
X63 25 20 18 GND n_mos $T=180100 -1810 0 0 $X=178900 $Y=-7090
X64 25 21 A2 GND n_mos $T=202200 27380 0 0 $X=201000 $Y=22100
X65 21 24 B2 GND n_mos $T=219580 27380 0 0 $X=218380 $Y=22100
X66 31 28 C2 GND n_mos $T=296160 -1810 0 0 $X=294960 $Y=-7090
X67 31 30 A3 GND n_mos $T=316660 27380 0 0 $X=315460 $Y=22100
X68 38 33 31 GND n_mos $T=347970 -1810 0 0 $X=346770 $Y=-7090
X69 38 34 A3 GND n_mos $T=370070 27380 0 0 $X=368870 $Y=22100
X70 34 37 B3 GND n_mos $T=387450 27380 0 0 $X=386250 $Y=22100
X71 44 41 C3 GND n_mos $T=466310 -1810 0 0 $X=465110 $Y=-7090
X72 44 43 A4 GND n_mos $T=486810 27380 0 0 $X=485610 $Y=22100
X73 51 46 44 GND n_mos $T=518120 -1810 0 0 $X=516920 $Y=-7090
X74 51 47 A4 GND n_mos $T=540220 27380 0 0 $X=539020 $Y=22100
X75 47 50 B4 GND n_mos $T=557600 27380 0 0 $X=556400 $Y=22100
X76 1 A1 VDD p_mos_VDD $T=-69430 8470 0 0 $X=-70630 $Y=7860
X77 1 B1 VDD p_mos_VDD $T=-55100 8470 0 0 $X=-56300 $Y=7860
X78 3 A1 VDD p_mos_VDD $T=-20080 34270 0 0 $X=-21280 $Y=33660
X79 9 A1 VDD p_mos_VDD $T=-5730 8030 0 0 $X=-6930 $Y=7420
X80 9 B1 VDD p_mos_VDD $T=32660 8030 0 0 $X=31460 $Y=7420
X81 6 A1 VDD p_mos_VDD $T=33580 34270 0 0 $X=32380 $Y=33660
X82 9 Cin VDD p_mos_VDD $T=45910 8030 0 0 $X=44710 $Y=7420
X83 14 A2 VDD p_mos_VDD $T=99200 8470 0 0 $X=98000 $Y=7860
X84 14 B2 VDD p_mos_VDD $T=113530 8470 0 0 $X=112330 $Y=7860
X85 16 A2 VDD p_mos_VDD $T=148550 34270 0 0 $X=147350 $Y=33660
X86 22 A2 VDD p_mos_VDD $T=162900 8030 0 0 $X=161700 $Y=7420
X87 22 B2 VDD p_mos_VDD $T=201290 8030 0 0 $X=200090 $Y=7420
X88 19 A2 VDD p_mos_VDD $T=202210 34270 0 0 $X=201010 $Y=33660
X89 22 C1 VDD p_mos_VDD $T=214540 8030 0 0 $X=213340 $Y=7420
X90 27 A3 VDD p_mos_VDD $T=267070 8470 0 0 $X=265870 $Y=7860
X91 27 B3 VDD p_mos_VDD $T=281400 8470 0 0 $X=280200 $Y=7860
X92 29 A3 VDD p_mos_VDD $T=316420 34270 0 0 $X=315220 $Y=33660
X93 35 A3 VDD p_mos_VDD $T=330770 8030 0 0 $X=329570 $Y=7420
X94 35 B3 VDD p_mos_VDD $T=369160 8030 0 0 $X=367960 $Y=7420
X95 32 A3 VDD p_mos_VDD $T=370080 34270 0 0 $X=368880 $Y=33660
X96 35 C2 VDD p_mos_VDD $T=382410 8030 0 0 $X=381210 $Y=7420
X97 40 A4 VDD p_mos_VDD $T=437220 8470 0 0 $X=436020 $Y=7860
X98 40 B4 VDD p_mos_VDD $T=451550 8470 0 0 $X=450350 $Y=7860
X99 42 A4 VDD p_mos_VDD $T=486570 34270 0 0 $X=485370 $Y=33660
X100 48 A4 VDD p_mos_VDD $T=500920 8030 0 0 $X=499720 $Y=7420
X101 48 B4 VDD p_mos_VDD $T=539310 8030 0 0 $X=538110 $Y=7420
X102 45 A4 VDD p_mos_VDD $T=540230 34270 0 0 $X=539030 $Y=33660
X103 48 C3 VDD p_mos_VDD $T=552560 8030 0 0 $X=551360 $Y=7420
.ENDS
***************************************
